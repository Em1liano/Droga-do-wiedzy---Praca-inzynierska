    ����          FAssembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null   
PlayerData   NameposXposYposZlevel
experiencedamagehealthmanacurrentQuestcurrentWorld         Quest         elo320(_bB Y;=TFC          B�     �C
   