    ����          FAssembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null   
PlayerData   NameposXposYposZlevel
experiencedamagehealthmanacurrentQuestcurrentWorld         Quest         	siemaEniuJ*�B��<p�}C          B�     �C	         Quest   isActivetitledescriptionexperienceRewardgoal  	QuestGoal       

    	      	QuestGoal   goalTyperequiredAmountcurrentAmount  GoalType      ����GoalType   value__                