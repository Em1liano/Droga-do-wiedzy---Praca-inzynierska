    ����          FAssembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null   
PlayerData   NameposXposYposZlevel
experiencedamagehealthmanacurrentQuestcurrentWorld         Quest         Emiliano�2p�<} C          B�     �C
   